`timescale 1ns/1ps 

module Timer_counter(
	input wire clk, reset, Start, Initial,
	output logic Ovf5);
	
	

endmodule